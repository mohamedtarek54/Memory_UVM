package memory_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "my_sequence_item.sv"
`include "my_sequence.sv"

`include "my_driver.sv"
`include "my_monitor.sv"
`include "my_sequencer.sv"
`include "my_agent.sv"
`include "my_scoreboard.sv"
`include "my_subscriber.sv"

`include "my_env.sv"

`include "my_test.sv"

endpackage : memory_pkg